library verilog;
use verilog.vl_types.all;
entity rle_testbench is
end rle_testbench;
