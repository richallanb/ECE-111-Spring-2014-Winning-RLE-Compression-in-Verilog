library verilog;
use verilog.vl_types.all;
entity tester is
end tester;
