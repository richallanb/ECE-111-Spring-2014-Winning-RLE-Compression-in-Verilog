library verilog;
use verilog.vl_types.all;
entity rle_testbench2 is
end rle_testbench2;
